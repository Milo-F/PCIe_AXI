`timescale 1ns/1ps
module tb_tlp_demux();
    
endmodule